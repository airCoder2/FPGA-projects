module lcd_controler (
    input clock, 
    output reg [0..7] DATA, LCD_EN, LCD_ON, LCD_RS, LCD_RW   
);





endmodule